magic
tech sky130A
magscale 1 2
timestamp 1717010029
<< pwell >>
rect 9528 274 9596 394
rect 12272 -1198 12340 -1100
<< viali >>
rect 7220 724 7610 768
rect 8036 258 8080 1032
rect 10682 272 10728 1028
rect 11134 734 11178 1004
rect 12420 734 12468 1004
rect 13684 738 13730 1032
rect 14208 726 14596 768
rect 8038 -1036 8082 -260
rect 8926 -1036 8968 -260
rect 12794 -558 12840 216
rect 13680 -558 13726 216
rect 8036 -1850 8080 -1556
rect 8922 -1850 8966 -1556
rect 9322 -1852 9374 -1582
rect 10612 -1852 10660 -1582
rect 11132 -1854 11176 -1098
rect 12796 -1852 12842 -1078
rect 13684 -1852 13726 -1078
<< metal1 >>
rect 7096 1396 14726 1502
rect 8036 1140 8084 1396
rect 12326 1232 12938 1270
rect 8024 1032 8094 1140
rect 7104 768 7726 788
rect 7104 724 7220 768
rect 7610 724 7726 768
rect 7104 712 7726 724
rect 7236 576 7296 664
rect 8024 258 8036 1032
rect 8080 670 8094 1032
rect 10674 1028 10744 1144
rect 10674 888 10682 1028
rect 10594 826 10682 888
rect 8080 624 8186 670
rect 8830 630 9534 682
rect 8080 258 8094 624
rect 8024 -260 8094 258
rect 8024 -1036 8038 -260
rect 8082 -630 8094 -260
rect 8460 -282 8520 294
rect 9528 274 9596 394
rect 10452 34 10520 302
rect 10674 272 10682 826
rect 10728 888 10744 1028
rect 11122 1004 11192 1116
rect 11122 888 11134 1004
rect 10728 826 11134 888
rect 10728 272 10744 826
rect 11122 734 11134 826
rect 11178 888 11192 1004
rect 12326 908 12370 1232
rect 12408 1004 12484 1118
rect 11178 826 11266 888
rect 11178 734 11192 826
rect 11122 624 11192 734
rect 10674 164 10744 272
rect 11340 34 11412 786
rect 12408 734 12420 1004
rect 12468 734 12484 1004
rect 12894 908 12938 1232
rect 13690 1144 13738 1396
rect 13672 1032 13746 1144
rect 13672 898 13684 1032
rect 12958 836 12960 888
rect 13584 856 13684 898
rect 12408 622 12484 734
rect 10452 -40 11412 34
rect 10452 -42 10520 -40
rect 8914 -260 8978 -142
rect 8786 -396 8852 -264
rect 8082 -674 8182 -630
rect 8082 -1036 8094 -674
rect 8024 -1142 8094 -1036
rect 8460 -1294 8520 -1012
rect 7574 -1346 8520 -1294
rect 7218 -2198 7258 -1388
rect 8024 -1556 8094 -1450
rect 8024 -1850 8036 -1556
rect 8080 -1682 8094 -1556
rect 8460 -1588 8520 -1346
rect 8914 -1036 8926 -260
rect 8968 -1036 8978 -260
rect 12418 -380 12472 622
rect 8914 -1556 8978 -1036
rect 9316 -448 12472 -380
rect 12784 216 12856 332
rect 9316 -1470 9380 -448
rect 12784 -558 12794 216
rect 12840 -558 12856 216
rect 13202 198 13262 774
rect 13672 738 13684 856
rect 13730 738 13746 1032
rect 13672 216 13746 738
rect 14100 768 14710 782
rect 14100 726 14208 768
rect 14596 726 14710 768
rect 14100 714 14710 726
rect 14522 570 14582 658
rect 13672 -156 13680 216
rect 13580 -196 13680 -156
rect 12916 -548 12982 -416
rect 10440 -856 11400 -782
rect 8080 -1724 8176 -1682
rect 8080 -1850 8094 -1724
rect 8024 -1954 8094 -1850
rect 8826 -2016 8874 -1702
rect 8914 -1850 8922 -1556
rect 8966 -1850 8978 -1556
rect 8914 -1964 8978 -1850
rect 9306 -1582 9384 -1470
rect 9306 -1852 9322 -1582
rect 9374 -1852 9384 -1582
rect 10440 -1608 10512 -856
rect 11120 -1098 11184 -980
rect 10604 -1582 10678 -1470
rect 10604 -1680 10612 -1582
rect 9306 -1962 9384 -1852
rect 9416 -2016 9464 -1702
rect 10522 -1742 10612 -1680
rect 10604 -1852 10612 -1742
rect 10660 -1680 10678 -1582
rect 11120 -1680 11132 -1098
rect 10660 -1742 11132 -1680
rect 10660 -1852 10678 -1742
rect 10604 -1964 10678 -1852
rect 8826 -2068 9464 -2016
rect 10824 -2198 10916 -1742
rect 11120 -1854 11132 -1742
rect 11176 -1680 11184 -1098
rect 11332 -1126 11400 -856
rect 12784 -1078 12856 -558
rect 12272 -1198 12340 -1100
rect 11176 -1742 11270 -1680
rect 11176 -1854 11184 -1742
rect 11120 -1962 11184 -1854
rect 12340 -2020 12384 -1726
rect 12784 -1852 12796 -1078
rect 12842 -1852 12856 -1078
rect 13272 -812 13332 -526
rect 13672 -558 13680 -196
rect 13726 -558 13746 216
rect 13672 -672 13746 -558
rect 13272 -864 14250 -812
rect 13272 -1102 13332 -864
rect 13674 -1078 13742 -966
rect 13674 -1446 13684 -1078
rect 13582 -1486 13684 -1446
rect 12784 -1964 12856 -1852
rect 12892 -2020 12936 -1726
rect 13674 -1852 13684 -1486
rect 13726 -1852 13742 -1078
rect 13674 -1966 13742 -1852
rect 12340 -2072 12936 -2020
rect 14562 -2198 14602 -1386
rect 7096 -2304 14726 -2198
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_0 ~/Desktop/MNEL
timestamp 1713891343
transform 1 0 11800 0 1 869
box -696 -267 696 267
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_1
timestamp 1713891343
transform 1 0 9992 0 1 -1717
box -696 -267 696 267
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_0 ~/Desktop/MNEL
timestamp 1713891343
transform 1 0 11796 0 1 -1476
box -696 -510 696 510
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_1
timestamp 1713891343
transform 1 0 10062 0 1 650
box -696 -510 696 510
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_0 ~/Desktop/MNEL
timestamp 1713898952
transform 1 0 7414 0 1 -419
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_1
timestamp 1713898952
transform 1 0 14402 0 1 -419
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_0 ~/Desktop/MNEL
timestamp 1713888985
transform 1 0 13264 0 1 885
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_1
timestamp 1713888985
transform 1 0 8500 0 1 -1703
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_0 ~/Desktop/MNEL
timestamp 1713888985
transform -1 0 8503 0 -1 -648
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_1
timestamp 1713888985
transform -1 0 13262 0 -1 -1465
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_2
timestamp 1713888985
transform -1 0 8502 0 -1 645
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_3
timestamp 1713888985
transform -1 0 13260 0 -1 -171
box -496 -519 496 519
<< end >>
