VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Saitama224_comp
  CLASS BLOCK ;
  FOREIGN tt_um_Saitama224_comp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 111.890 16.830 115.150 29.020 ;
        RECT 116.480 25.650 121.440 30.840 ;
      LAYER pwell ;
        RECT 123.280 25.720 130.240 30.820 ;
        RECT 131.970 28.030 138.930 30.700 ;
      LAYER nwell ;
        RECT 140.290 28.050 145.250 30.840 ;
        RECT 116.485 19.185 121.445 24.375 ;
        RECT 140.270 21.570 145.230 26.760 ;
        RECT 116.470 15.110 121.430 17.900 ;
      LAYER pwell ;
        RECT 122.930 15.100 129.890 17.770 ;
        RECT 131.950 15.090 138.910 20.190 ;
      LAYER nwell ;
        RECT 140.280 15.100 145.240 20.290 ;
        RECT 146.830 16.830 150.090 29.020 ;
      LAYER li1 ;
        RECT 116.660 30.490 121.260 30.660 ;
        RECT 116.660 30.180 116.830 30.490 ;
        RECT 112.550 28.840 114.500 28.860 ;
        RECT 112.070 28.670 114.970 28.840 ;
        RECT 112.070 17.180 112.240 28.670 ;
        RECT 112.550 28.640 114.500 28.670 ;
        RECT 112.870 28.160 114.170 28.330 ;
        RECT 112.640 17.905 112.810 27.945 ;
        RECT 114.230 17.905 114.400 27.945 ;
        RECT 112.870 17.520 114.170 17.690 ;
        RECT 114.800 17.180 114.970 28.670 ;
        RECT 116.630 26.310 116.850 30.180 ;
        RECT 117.460 29.980 120.460 30.150 ;
        RECT 117.230 26.725 117.400 29.765 ;
        RECT 120.520 26.725 120.690 29.765 ;
        RECT 117.460 26.340 120.460 26.510 ;
        RECT 116.660 26.000 116.830 26.310 ;
        RECT 121.090 26.000 121.260 30.490 ;
        RECT 116.660 25.830 121.260 26.000 ;
        RECT 123.460 30.470 130.060 30.640 ;
        RECT 123.460 26.070 123.630 30.470 ;
        RECT 129.890 30.160 130.060 30.470 ;
        RECT 132.150 30.350 138.750 30.520 ;
        RECT 124.260 29.960 129.260 30.130 ;
        RECT 124.030 26.750 124.200 29.790 ;
        RECT 129.320 26.750 129.490 29.790 ;
        RECT 124.260 26.410 129.260 26.580 ;
        RECT 129.860 26.380 130.090 30.160 ;
        RECT 132.150 30.040 132.320 30.350 ;
        RECT 138.580 30.040 138.750 30.350 ;
        RECT 140.470 30.490 145.070 30.660 ;
        RECT 132.120 28.690 132.340 30.040 ;
        RECT 132.950 29.840 137.950 30.010 ;
        RECT 132.720 29.060 132.890 29.670 ;
        RECT 138.010 29.060 138.180 29.670 ;
        RECT 132.950 28.720 137.950 28.890 ;
        RECT 138.550 28.690 138.790 30.040 ;
        RECT 132.150 28.380 132.320 28.690 ;
        RECT 138.580 28.380 138.750 28.690 ;
        RECT 132.150 28.210 138.750 28.380 ;
        RECT 140.470 28.400 140.640 30.490 ;
        RECT 144.900 30.180 145.070 30.490 ;
        RECT 141.270 29.980 144.270 30.150 ;
        RECT 141.040 29.125 141.210 29.765 ;
        RECT 144.330 29.125 144.500 29.765 ;
        RECT 141.270 28.740 144.270 28.910 ;
        RECT 144.870 28.710 145.100 30.180 ;
        RECT 147.490 28.840 149.430 28.860 ;
        RECT 144.900 28.400 145.070 28.710 ;
        RECT 140.470 28.230 145.070 28.400 ;
        RECT 147.010 28.670 149.910 28.840 ;
        RECT 140.450 26.410 145.050 26.580 ;
        RECT 129.890 26.070 130.060 26.380 ;
        RECT 140.450 26.100 140.620 26.410 ;
        RECT 144.880 26.100 145.050 26.410 ;
        RECT 123.460 25.900 130.060 26.070 ;
        RECT 116.665 24.025 121.265 24.195 ;
        RECT 116.665 23.720 116.835 24.025 ;
        RECT 121.095 23.720 121.265 24.025 ;
        RECT 116.640 19.840 116.860 23.720 ;
        RECT 117.465 23.515 120.465 23.685 ;
        RECT 117.235 20.260 117.405 23.300 ;
        RECT 120.525 20.260 120.695 23.300 ;
        RECT 117.465 19.875 120.465 20.045 ;
        RECT 121.080 19.840 121.290 23.720 ;
        RECT 140.420 22.230 140.650 26.100 ;
        RECT 141.250 25.900 144.250 26.070 ;
        RECT 141.020 22.645 141.190 25.685 ;
        RECT 144.310 22.645 144.480 25.685 ;
        RECT 141.250 22.260 144.250 22.430 ;
        RECT 144.850 22.230 145.080 26.100 ;
        RECT 140.450 21.920 140.620 22.230 ;
        RECT 144.880 21.920 145.050 22.230 ;
        RECT 140.450 21.750 145.050 21.920 ;
        RECT 132.130 19.840 138.730 20.010 ;
        RECT 116.665 19.535 116.835 19.840 ;
        RECT 121.095 19.535 121.265 19.840 ;
        RECT 116.665 19.365 121.265 19.535 ;
        RECT 132.130 19.530 132.300 19.840 ;
        RECT 116.650 17.550 121.250 17.720 ;
        RECT 116.650 17.240 116.820 17.550 ;
        RECT 121.080 17.240 121.250 17.550 ;
        RECT 123.110 17.420 129.710 17.590 ;
        RECT 112.070 17.010 114.970 17.180 ;
        RECT 116.630 15.770 116.850 17.240 ;
        RECT 117.450 17.040 120.450 17.210 ;
        RECT 117.220 16.185 117.390 16.825 ;
        RECT 120.510 16.185 120.680 16.825 ;
        RECT 117.450 15.800 120.450 15.970 ;
        RECT 121.060 15.770 121.280 17.240 ;
        RECT 123.110 17.110 123.280 17.420 ;
        RECT 129.540 17.110 129.710 17.420 ;
        RECT 116.650 15.460 116.820 15.770 ;
        RECT 121.080 15.460 121.250 15.770 ;
        RECT 123.060 15.760 123.320 17.110 ;
        RECT 123.910 16.910 128.910 17.080 ;
        RECT 123.680 16.130 123.850 16.740 ;
        RECT 128.970 16.130 129.140 16.740 ;
        RECT 123.910 15.790 128.910 15.960 ;
        RECT 129.510 15.760 129.750 17.110 ;
        RECT 116.650 15.290 121.250 15.460 ;
        RECT 123.110 15.450 123.280 15.760 ;
        RECT 129.540 15.450 129.710 15.760 ;
        RECT 132.110 15.750 132.330 19.530 ;
        RECT 132.930 19.330 137.930 19.500 ;
        RECT 132.700 16.120 132.870 19.160 ;
        RECT 137.990 16.120 138.160 19.160 ;
        RECT 132.930 15.780 137.930 15.950 ;
        RECT 123.110 15.280 129.710 15.450 ;
        RECT 132.130 15.440 132.300 15.750 ;
        RECT 138.560 15.440 138.730 19.840 ;
        RECT 140.460 19.940 145.060 20.110 ;
        RECT 140.460 19.630 140.630 19.940 ;
        RECT 144.890 19.630 145.060 19.940 ;
        RECT 140.430 15.760 140.660 19.630 ;
        RECT 141.260 19.430 144.260 19.600 ;
        RECT 141.030 16.175 141.200 19.215 ;
        RECT 144.320 16.175 144.490 19.215 ;
        RECT 141.260 15.790 144.260 15.960 ;
        RECT 144.870 15.760 145.080 19.630 ;
        RECT 147.010 17.180 147.180 28.670 ;
        RECT 147.490 28.650 149.430 28.670 ;
        RECT 147.810 28.160 149.110 28.330 ;
        RECT 147.580 17.905 147.750 27.945 ;
        RECT 149.170 17.905 149.340 27.945 ;
        RECT 147.810 17.520 149.110 17.690 ;
        RECT 149.740 17.180 149.910 28.670 ;
        RECT 147.010 17.010 149.910 17.180 ;
        RECT 132.130 15.270 138.730 15.440 ;
        RECT 140.460 15.450 140.630 15.760 ;
        RECT 144.890 15.450 145.060 15.760 ;
        RECT 140.460 15.280 145.060 15.450 ;
      LAYER mcon ;
        RECT 112.950 28.160 114.090 28.330 ;
        RECT 112.640 17.985 112.810 27.865 ;
        RECT 114.230 17.985 114.400 27.865 ;
        RECT 112.950 17.520 114.090 17.690 ;
        RECT 116.630 26.310 116.850 30.180 ;
        RECT 117.540 29.980 120.380 30.150 ;
        RECT 117.230 26.805 117.400 29.685 ;
        RECT 120.520 26.805 120.690 29.685 ;
        RECT 117.540 26.340 120.380 26.510 ;
        RECT 124.340 29.960 129.180 30.130 ;
        RECT 124.030 26.830 124.200 29.710 ;
        RECT 129.320 26.830 129.490 29.710 ;
        RECT 124.340 26.410 129.180 26.580 ;
        RECT 129.860 26.380 130.090 30.160 ;
        RECT 132.120 28.690 132.340 30.040 ;
        RECT 133.030 29.840 137.870 30.010 ;
        RECT 132.720 29.140 132.890 29.590 ;
        RECT 138.010 29.140 138.180 29.590 ;
        RECT 133.030 28.720 137.870 28.890 ;
        RECT 138.550 28.690 138.790 30.040 ;
        RECT 141.350 29.980 144.190 30.150 ;
        RECT 141.040 29.205 141.210 29.685 ;
        RECT 144.330 29.205 144.500 29.685 ;
        RECT 141.350 28.740 144.190 28.910 ;
        RECT 144.870 28.710 145.100 30.180 ;
        RECT 117.545 23.515 120.385 23.685 ;
        RECT 117.235 20.340 117.405 23.220 ;
        RECT 120.525 20.340 120.695 23.220 ;
        RECT 117.545 19.875 120.385 20.045 ;
        RECT 140.420 22.230 140.650 26.100 ;
        RECT 141.330 25.900 144.170 26.070 ;
        RECT 141.020 22.725 141.190 25.605 ;
        RECT 144.310 22.725 144.480 25.605 ;
        RECT 141.330 22.260 144.170 22.430 ;
        RECT 144.850 22.230 145.080 26.100 ;
        RECT 116.630 15.770 116.850 17.240 ;
        RECT 117.530 17.040 120.370 17.210 ;
        RECT 117.220 16.265 117.390 16.745 ;
        RECT 120.510 16.265 120.680 16.745 ;
        RECT 117.530 15.800 120.370 15.970 ;
        RECT 121.060 15.770 121.280 17.240 ;
        RECT 123.060 15.760 123.320 17.110 ;
        RECT 123.990 16.910 128.830 17.080 ;
        RECT 123.680 16.210 123.850 16.660 ;
        RECT 128.970 16.210 129.140 16.660 ;
        RECT 123.990 15.790 128.830 15.960 ;
        RECT 129.510 15.760 129.750 17.110 ;
        RECT 132.110 15.750 132.330 19.530 ;
        RECT 133.010 19.330 137.850 19.500 ;
        RECT 132.700 16.200 132.870 19.080 ;
        RECT 137.990 16.200 138.160 19.080 ;
        RECT 133.010 15.780 137.850 15.950 ;
        RECT 140.430 15.760 140.660 19.630 ;
        RECT 141.340 19.430 144.180 19.600 ;
        RECT 141.030 16.255 141.200 19.135 ;
        RECT 144.320 16.255 144.490 19.135 ;
        RECT 141.340 15.790 144.180 15.960 ;
        RECT 144.870 15.760 145.080 19.630 ;
        RECT 147.890 28.160 149.030 28.330 ;
        RECT 147.580 17.985 147.750 27.865 ;
        RECT 149.170 17.985 149.340 27.865 ;
        RECT 147.890 17.520 149.030 17.690 ;
      LAYER met1 ;
        RECT 151.020 34.210 152.020 34.240 ;
        RECT 106.040 32.530 109.030 33.350 ;
        RECT 113.090 33.210 152.020 34.210 ;
        RECT 151.020 33.180 152.020 33.210 ;
        RECT 106.040 32.000 150.080 32.530 ;
        RECT 106.040 31.730 109.030 32.000 ;
        RECT 113.120 28.960 114.120 31.710 ;
        RECT 116.630 30.720 116.870 32.000 ;
        RECT 138.080 31.180 141.140 31.370 ;
        RECT 111.970 28.580 115.080 28.960 ;
        RECT 116.570 28.370 116.920 30.720 ;
        RECT 117.480 29.950 120.440 30.180 ;
        RECT 124.280 29.930 129.240 30.160 ;
        RECT 117.200 28.370 117.430 29.745 ;
        RECT 112.890 28.340 114.150 28.360 ;
        RECT 112.630 28.130 114.150 28.340 ;
        RECT 116.570 28.140 117.430 28.370 ;
        RECT 112.630 27.925 112.930 28.130 ;
        RECT 112.610 27.900 112.930 27.925 ;
        RECT 112.610 18.080 112.840 27.900 ;
        RECT 112.540 17.925 112.840 18.080 ;
        RECT 114.200 18.550 114.430 27.925 ;
        RECT 116.570 21.870 116.920 28.140 ;
        RECT 117.200 26.745 117.430 28.140 ;
        RECT 120.490 28.430 120.720 29.745 ;
        RECT 124.000 28.430 124.230 29.770 ;
        RECT 120.490 28.170 124.230 28.430 ;
        RECT 120.490 26.745 120.720 28.170 ;
        RECT 124.000 26.990 124.230 28.170 ;
        RECT 129.290 29.460 129.520 29.770 ;
        RECT 129.820 29.460 130.170 30.740 ;
        RECT 132.060 29.460 132.410 30.600 ;
        RECT 132.970 29.810 137.930 30.040 ;
        RECT 138.080 29.650 138.300 31.180 ;
        RECT 132.690 29.460 132.920 29.650 ;
        RECT 129.290 29.150 132.920 29.460 ;
        RECT 124.000 26.770 124.430 26.990 ;
        RECT 129.290 26.770 129.520 29.150 ;
        RECT 124.090 26.610 124.430 26.770 ;
        RECT 117.480 26.310 120.440 26.540 ;
        RECT 124.090 26.390 129.240 26.610 ;
        RECT 124.280 26.380 129.240 26.390 ;
        RECT 118.750 23.715 119.050 26.310 ;
        RECT 128.710 25.190 129.050 26.380 ;
        RECT 129.820 25.840 130.170 29.150 ;
        RECT 132.060 28.140 132.410 29.150 ;
        RECT 132.690 29.080 132.920 29.150 ;
        RECT 137.980 29.560 138.300 29.650 ;
        RECT 137.980 29.080 138.210 29.560 ;
        RECT 133.150 28.920 133.510 28.950 ;
        RECT 132.970 28.690 137.930 28.920 ;
        RECT 133.150 25.190 133.510 28.690 ;
        RECT 138.490 28.130 138.870 30.610 ;
        RECT 140.920 29.745 141.140 31.180 ;
        RECT 144.900 30.740 145.140 32.000 ;
        RECT 150.700 30.810 151.700 30.840 ;
        RECT 141.290 29.950 144.250 30.180 ;
        RECT 140.920 29.560 141.240 29.745 ;
        RECT 141.010 29.460 141.240 29.560 ;
        RECT 144.300 29.510 144.530 29.745 ;
        RECT 144.810 29.510 145.180 30.740 ;
        RECT 148.365 29.810 151.700 30.810 ;
        RECT 141.010 29.200 141.250 29.460 ;
        RECT 144.300 29.300 145.180 29.510 ;
        RECT 141.010 29.145 141.240 29.200 ;
        RECT 144.300 29.145 144.530 29.300 ;
        RECT 141.290 28.710 144.250 28.940 ;
        RECT 128.710 24.820 133.510 25.190 ;
        RECT 128.710 24.810 129.050 24.820 ;
        RECT 117.485 23.700 120.445 23.715 ;
        RECT 117.485 23.485 120.710 23.700 ;
        RECT 120.380 23.280 120.710 23.485 ;
        RECT 117.205 21.870 117.435 23.280 ;
        RECT 120.380 23.040 120.725 23.280 ;
        RECT 116.570 21.650 117.435 21.870 ;
        RECT 116.570 19.310 116.920 21.650 ;
        RECT 117.205 20.280 117.435 21.650 ;
        RECT 120.495 20.280 120.725 23.040 ;
        RECT 117.485 19.845 120.445 20.075 ;
        RECT 118.750 18.550 119.050 19.845 ;
        RECT 114.200 18.290 119.050 18.550 ;
        RECT 114.200 17.925 114.430 18.290 ;
        RECT 104.000 14.030 109.020 14.830 ;
        RECT 112.540 14.030 112.740 17.925 ;
        RECT 112.890 17.490 114.150 17.720 ;
        RECT 116.570 16.610 116.920 17.770 ;
        RECT 118.750 17.240 119.050 18.290 ;
        RECT 117.470 17.010 120.430 17.240 ;
        RECT 117.190 16.610 117.420 16.805 ;
        RECT 116.570 16.400 117.420 16.610 ;
        RECT 116.570 15.250 116.920 16.400 ;
        RECT 117.190 16.205 117.420 16.400 ;
        RECT 120.480 16.510 120.710 16.805 ;
        RECT 120.480 16.205 120.820 16.510 ;
        RECT 117.470 15.770 120.430 16.000 ;
        RECT 120.580 14.940 120.820 16.205 ;
        RECT 121.020 15.200 121.340 24.310 ;
        RECT 138.540 23.120 138.810 28.130 ;
        RECT 123.030 22.780 138.810 23.120 ;
        RECT 123.030 17.670 123.350 22.780 ;
        RECT 128.650 20.740 133.450 21.110 ;
        RECT 122.980 15.210 123.370 17.670 ;
        RECT 128.650 17.110 129.010 20.740 ;
        RECT 123.930 16.980 129.010 17.110 ;
        RECT 123.930 16.880 128.890 16.980 ;
        RECT 123.650 16.510 123.880 16.720 ;
        RECT 123.530 16.150 123.880 16.510 ;
        RECT 128.940 16.620 129.170 16.720 ;
        RECT 129.470 16.620 129.840 17.670 ;
        RECT 132.050 16.620 132.370 20.120 ;
        RECT 133.110 19.530 133.450 20.740 ;
        RECT 132.950 19.520 137.910 19.530 ;
        RECT 132.950 19.300 138.150 19.520 ;
        RECT 137.810 19.140 138.150 19.300 ;
        RECT 132.670 16.620 132.900 19.140 ;
        RECT 137.810 19.030 138.190 19.140 ;
        RECT 128.940 16.310 132.900 16.620 ;
        RECT 128.940 16.150 129.170 16.310 ;
        RECT 121.700 14.940 122.660 15.210 ;
        RECT 123.530 14.940 123.770 16.150 ;
        RECT 123.930 15.760 128.890 15.990 ;
        RECT 129.470 15.200 129.840 16.310 ;
        RECT 120.580 14.680 123.770 14.940 ;
        RECT 121.700 14.250 122.660 14.680 ;
        RECT 130.570 14.030 131.030 16.310 ;
        RECT 132.050 15.210 132.370 16.310 ;
        RECT 132.670 16.140 132.900 16.310 ;
        RECT 137.960 16.390 138.190 19.030 ;
        RECT 137.960 16.140 138.370 16.390 ;
        RECT 132.950 15.750 137.910 15.980 ;
        RECT 138.150 14.920 138.370 16.140 ;
        RECT 140.370 15.200 140.730 26.680 ;
        RECT 142.460 26.100 142.760 28.710 ;
        RECT 141.270 25.870 144.230 26.100 ;
        RECT 140.990 22.940 141.220 25.665 ;
        RECT 144.280 24.240 144.510 25.665 ;
        RECT 144.810 24.240 145.180 29.300 ;
        RECT 148.385 28.930 149.350 29.810 ;
        RECT 150.700 29.780 151.700 29.810 ;
        RECT 146.950 28.590 150.000 28.930 ;
        RECT 147.830 28.310 149.090 28.360 ;
        RECT 147.830 28.130 149.360 28.310 ;
        RECT 149.060 27.925 149.360 28.130 ;
        RECT 144.280 24.040 145.180 24.240 ;
        RECT 140.990 22.665 141.360 22.940 ;
        RECT 144.280 22.665 144.510 24.040 ;
        RECT 141.030 22.460 141.360 22.665 ;
        RECT 141.030 22.280 144.230 22.460 ;
        RECT 141.270 22.230 144.230 22.280 ;
        RECT 142.810 20.960 143.110 22.230 ;
        RECT 144.810 21.660 145.180 24.040 ;
        RECT 147.550 20.960 147.780 27.925 ;
        RECT 149.060 27.870 149.370 27.925 ;
        RECT 142.810 20.700 147.780 20.960 ;
        RECT 142.810 19.630 143.110 20.700 ;
        RECT 141.280 19.400 144.240 19.630 ;
        RECT 141.000 16.390 141.230 19.195 ;
        RECT 140.910 16.195 141.230 16.390 ;
        RECT 144.290 17.790 144.520 19.195 ;
        RECT 144.820 17.790 145.160 20.190 ;
        RECT 147.550 17.925 147.780 20.700 ;
        RECT 149.140 18.090 149.370 27.870 ;
        RECT 149.140 17.925 149.460 18.090 ;
        RECT 144.290 17.590 145.160 17.790 ;
        RECT 144.290 16.195 144.520 17.590 ;
        RECT 140.910 14.920 141.130 16.195 ;
        RECT 141.280 15.760 144.240 15.990 ;
        RECT 144.820 15.190 145.160 17.590 ;
        RECT 147.830 17.490 149.090 17.720 ;
        RECT 138.150 14.660 141.130 14.920 ;
        RECT 149.260 14.030 149.460 17.925 ;
        RECT 104.000 13.500 150.080 14.030 ;
        RECT 104.000 13.210 109.020 13.500 ;
      LAYER via ;
        RECT 106.080 31.730 107.700 33.350 ;
        RECT 113.120 33.210 114.120 34.210 ;
        RECT 151.020 33.210 152.020 34.210 ;
        RECT 113.120 30.680 114.120 31.680 ;
        RECT 150.700 29.810 151.700 30.810 ;
        RECT 104.040 13.210 105.660 14.830 ;
        RECT 121.730 14.280 122.630 15.180 ;
      LAYER met2 ;
        RECT 102.990 31.730 107.730 33.350 ;
        RECT 113.120 30.650 114.120 34.240 ;
        RECT 150.990 34.190 152.050 34.210 ;
        RECT 150.990 33.230 153.790 34.190 ;
        RECT 150.990 33.210 152.050 33.230 ;
        RECT 150.670 30.790 151.730 30.810 ;
        RECT 150.670 29.830 153.470 30.790 ;
        RECT 150.670 29.810 151.730 29.830 ;
        RECT 100.950 13.210 105.690 14.830 ;
        RECT 121.730 12.280 122.630 15.210 ;
      LAYER via2 ;
        RECT 103.040 31.770 104.580 33.310 ;
        RECT 152.780 33.230 153.740 34.190 ;
        RECT 152.460 29.830 153.420 30.790 ;
        RECT 101.000 13.250 102.540 14.790 ;
        RECT 121.755 12.325 122.605 13.175 ;
      LAYER met3 ;
        RECT 152.755 34.170 153.765 34.215 ;
        RECT 37.285 33.320 38.835 33.345 ;
        RECT 37.280 31.760 61.280 33.320 ;
        RECT 103.015 33.310 104.605 33.335 ;
        RECT 99.400 31.770 104.605 33.310 ;
        RECT 152.755 33.250 155.690 34.170 ;
        RECT 152.755 33.205 153.765 33.250 ;
        RECT 37.285 31.735 38.835 31.760 ;
        RECT 103.015 31.745 104.605 31.770 ;
        RECT 152.435 30.770 153.445 30.815 ;
        RECT 152.435 29.850 155.370 30.770 ;
        RECT 152.435 29.805 153.445 29.850 ;
        RECT 100.975 14.790 102.565 14.815 ;
        RECT 97.360 13.250 102.565 14.790 ;
        RECT 100.975 13.225 102.565 13.250 ;
        RECT 121.730 11.720 122.630 13.200 ;
        RECT 121.700 10.820 122.660 11.720 ;
      LAYER via3 ;
        RECT 37.285 31.765 38.835 33.315 ;
        RECT 59.695 31.765 61.245 33.315 ;
        RECT 99.435 31.775 100.965 33.305 ;
        RECT 154.740 33.250 155.660 34.170 ;
        RECT 154.420 29.850 155.340 30.770 ;
        RECT 97.395 13.255 98.925 14.785 ;
        RECT 121.730 10.820 122.630 11.720 ;
      LAYER met4 ;
        RECT 3.990 223.710 4.290 224.760 ;
        RECT 7.670 223.710 7.970 224.760 ;
        RECT 11.350 223.710 11.650 224.760 ;
        RECT 15.030 223.710 15.330 224.760 ;
        RECT 18.710 223.710 19.010 224.760 ;
        RECT 22.390 223.710 22.690 224.760 ;
        RECT 26.070 223.710 26.370 224.760 ;
        RECT 29.750 223.710 30.050 224.760 ;
        RECT 33.430 223.710 33.730 224.760 ;
        RECT 37.110 223.710 37.410 224.760 ;
        RECT 40.790 223.710 41.090 224.760 ;
        RECT 44.470 223.710 44.770 224.760 ;
        RECT 48.150 223.710 48.450 224.760 ;
        RECT 51.830 223.710 52.130 224.760 ;
        RECT 55.510 223.710 55.810 224.760 ;
        RECT 59.190 223.710 59.490 224.760 ;
        RECT 62.870 223.710 63.170 224.760 ;
        RECT 66.550 223.710 66.850 224.760 ;
        RECT 70.230 223.710 70.530 224.760 ;
        RECT 73.910 223.710 74.210 224.760 ;
        RECT 77.590 223.710 77.890 224.760 ;
        RECT 81.270 223.710 81.570 224.760 ;
        RECT 84.950 223.710 85.250 224.760 ;
        RECT 88.630 223.710 88.930 224.760 ;
        RECT 3.990 223.410 88.930 223.710 ;
        RECT 49.000 220.760 50.500 223.410 ;
        RECT 154.735 34.160 155.665 34.175 ;
        RECT 37.280 33.290 38.840 33.320 ;
        RECT 2.500 31.790 38.840 33.290 ;
        RECT 37.280 31.760 38.840 31.790 ;
        RECT 59.690 33.290 61.250 33.320 ;
        RECT 99.430 33.290 100.970 33.310 ;
        RECT 59.690 31.790 100.970 33.290 ;
        RECT 154.735 33.260 157.310 34.160 ;
        RECT 154.735 33.245 155.665 33.260 ;
        RECT 59.690 31.760 61.250 31.790 ;
        RECT 99.430 31.770 100.970 31.790 ;
        RECT 154.415 30.760 155.345 30.775 ;
        RECT 154.415 29.860 155.370 30.760 ;
        RECT 154.415 29.845 155.345 29.860 ;
        RECT 97.390 14.770 98.930 14.790 ;
        RECT 50.500 13.270 98.930 14.770 ;
        RECT 97.390 13.250 98.930 13.270 ;
        RECT 121.725 10.815 122.635 11.725 ;
        RECT 121.730 9.580 122.630 10.815 ;
        RECT 112.250 8.680 122.630 9.580 ;
        RECT 154.430 9.530 155.330 29.845 ;
        RECT 112.250 1.000 113.150 8.680 ;
        RECT 134.330 8.630 155.330 9.530 ;
        RECT 134.330 1.000 135.230 8.630 ;
        RECT 156.410 1.000 157.310 33.260 ;
  END
END tt_um_Saitama224_comp
END LIBRARY

